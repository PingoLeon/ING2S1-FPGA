-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition
-- Created on Thu Nov 02 17:30:57 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY porte IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        SW9 : IN STD_LOGIC := '0';
        SW8 : IN STD_LOGIC := '0';
        Pause : IN STD_LOGIC := '0';
        HEX15 : OUT STD_LOGIC;
        HEX24 : OUT STD_LOGIC;
        HEX3 : OUT STD_LOGIC
    );
END porte;

ARCHITECTURE BEHAVIOR OF porte IS
    TYPE type_fstate IS (ferme,moitie1,ouvert,moitie2);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,SW9,SW8,Pause)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= ferme;
            HEX15 <= '0';
            HEX24 <= '0';
            HEX3 <= '0';
        ELSE
            HEX15 <= '0';
            HEX24 <= '0';
            HEX3 <= '0';
            CASE fstate IS
                WHEN ferme =>
                    IF ((SW9 = '1')) THEN
                        reg_fstate <= moitie1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ferme;
                    END IF;

                    HEX3 <= '1';

                    HEX15 <= '1';

                    HEX24 <= '1';
                WHEN moitie1 =>
                    IF ((SW9 = '1')) THEN
                        reg_fstate <= moitie2;
                    ELSIF ((((SW8 = '1') AND NOT((SW9 = '1'))) AND NOT((Pause = '1')))) THEN
                        reg_fstate <= ferme;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= moitie1;
                    END IF;

                    HEX3 <= '0';

                    HEX15 <= '1';

                    HEX24 <= '1';
                WHEN ouvert =>
                    IF ((((SW8 = '1') AND NOT((SW9 = '1'))) AND NOT((Pause = '1')))) THEN
                        reg_fstate <= moitie2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= ouvert;
                    END IF;

                    HEX3 <= '0';

                    HEX15 <= '0';

                    HEX24 <= '0';
                WHEN moitie2 =>
                    IF ((SW9 = '1')) THEN
                        reg_fstate <= ouvert;
                    ELSIF ((((SW8 = '1') AND NOT((SW9 = '1'))) AND NOT((Pause = '1')))) THEN
                        reg_fstate <= moitie1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= moitie2;
                    END IF;

                    HEX3 <= '0';

                    HEX15 <= '1';

                    HEX24 <= '0';
                WHEN OTHERS => 
                    HEX15 <= 'X';
                    HEX24 <= 'X';
                    HEX3 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
