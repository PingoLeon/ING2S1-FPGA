-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition
-- Created on Thu Nov 02 13:32:30 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY MSMdpsmf IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        KEY0 : IN STD_LOGIC := '0';
        KEY1 : IN STD_LOGIC := '0';
        SW7 : IN STD_LOGIC := '0';
        CLK5 : IN STD_LOGIC := '0';
        MDP : OUT STD_LOGIC
    );
END MSMdpsmf;

ARCHITECTURE BEHAVIOR OF MSMdpsmf IS
    TYPE type_fstate IS (Init,state2,state3,state4,state5,state9,state,state6,state10,state7,state8);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_MDP : STD_LOGIC := '0';
BEGIN
    PROCESS (clock,reg_fstate,reg_MDP)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
            MDP <= reg_MDP;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,KEY0,KEY1,SW7,CLK5)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Init;
            reg_MDP <= '0';
        ELSE
            reg_MDP <= '0';
            CASE fstate IS
                WHEN Init =>
                    IF (((KEY0 = '1') AND (SW7 = '1'))) THEN
                        reg_fstate <= state;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Init;
                    END IF;

                    reg_MDP <= '0';
                WHEN state2 =>
                    IF ((((KEY0 = '1') AND (SW7 = '1')) AND NOT((CLK5 = '1')))) THEN
                        reg_fstate <= state3;
                    ELSIF ((CLK5 = '1')) THEN
                        reg_fstate <= Init;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    reg_MDP <= '0';
                WHEN state3 =>
                    IF ((NOT((KEY0 = '1')) AND (SW7 = '1'))) THEN
                        reg_fstate <= state4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    reg_MDP <= '0';
                WHEN state4 =>
                    IF ((((KEY1 = '1') AND (SW7 = '1')) AND NOT((CLK5 = '1')))) THEN
                        reg_fstate <= state5;
                    ELSIF ((CLK5 = '1')) THEN
                        reg_fstate <= Init;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state4;
                    END IF;

                    reg_MDP <= '0';
                WHEN state5 =>
                    IF ((NOT((KEY1 = '1')) AND (SW7 = '1'))) THEN
                        reg_fstate <= state6;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state5;
                    END IF;

                    reg_MDP <= '0';
                WHEN state9 =>
                    IF ((NOT((KEY0 = '1')) AND (SW7 = '1'))) THEN
                        reg_fstate <= state10;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state9;
                    END IF;

                    reg_MDP <= '0';
                WHEN state =>
                    IF ((NOT((KEY0 = '1')) AND (SW7 = '1'))) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state;
                    END IF;

                    reg_MDP <= '0';
                WHEN state6 =>
                    IF ((((KEY0 = '1') AND (SW7 = '1')) AND NOT((CLK5 = '1')))) THEN
                        reg_fstate <= state7;
                    ELSIF ((CLK5 = '1')) THEN
                        reg_fstate <= Init;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state6;
                    END IF;

                    reg_MDP <= '0';
                WHEN state10 =>
                    IF ((SW7 = '1')) THEN
                        reg_fstate <= state10;
                    ELSIF (NOT((SW7 = '1'))) THEN
                        reg_fstate <= Init;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state10;
                    END IF;

                    reg_MDP <= '1';
                WHEN state7 =>
                    IF ((NOT((KEY0 = '1')) AND (SW7 = '1'))) THEN
                        reg_fstate <= state8;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state7;
                    END IF;

                    reg_MDP <= '0';
                WHEN state8 =>
                    IF ((((KEY0 = '1') AND (SW7 = '1')) AND NOT((CLK5 = '1')))) THEN
                        reg_fstate <= state9;
                    ELSIF ((CLK5 = '1')) THEN
                        reg_fstate <= Init;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state8;
                    END IF;

                    reg_MDP <= '0';
                WHEN OTHERS => 
                    reg_MDP <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
