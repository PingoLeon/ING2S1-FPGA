-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition
-- Created on Fri Nov 03 12:32:57 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY cyclePorteFermee IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        SW1 : IN STD_LOGIC := '0';
        SW2 : IN STD_LOGIC := '0';
        SW3 : IN STD_LOGIC := '0';
        SW4 : IN STD_LOGIC := '0';
        SW5 : IN STD_LOGIC := '0';
        SW6 : IN STD_LOGIC := '0';
        SW7 : IN STD_LOGIC := '0';
        SW8 : IN STD_LOGIC := '0';
        E1 : IN STD_LOGIC := '0';
        E2 : IN STD_LOGIC := '0';
        E3 : IN STD_LOGIC := '0';
        E4 : IN STD_LOGIC := '0';
        E5 : IN STD_LOGIC := '0';
        E6 : IN STD_LOGIC := '0';
        E7 : IN STD_LOGIC := '0';
        E8 : IN STD_LOGIC := '0';
        Fermee : OUT STD_LOGIC
    );
END cyclePorteFermee;

ARCHITECTURE BEHAVIOR OF cyclePorteFermee IS
    TYPE type_fstate IS (state2,Base);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,SW1,SW2,SW3,SW4,SW5,SW6,SW7,SW8,E1,E2,E3,E4,E5,E6,E7,E8)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= Base;
            Fermee <= '0';
        ELSE
            Fermee <= '0';
            CASE fstate IS
                WHEN state2 =>
                    IF (NOT((((((((((E1 = '1') AND (SW1 = '1')) OR ((E2 = '1') AND (SW2 = '1'))) OR ((E3 = '1') AND (SW3 = '1'))) OR ((E4 = '1') AND (SW4 = '1'))) OR ((E5 = '1') AND (SW5 = '1'))) OR ((E6 = '1') AND (SW6 = '1'))) OR ((E7 = '1') AND (SW7 = '1'))) OR ((E8 = '1') AND (SW8 = '1'))))) THEN
                        reg_fstate <= Base;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    Fermee <= '0';
                WHEN Base =>
                    IF ((((((((((E1 = '1') AND (SW1 = '1')) OR ((E2 = '1') AND (SW2 = '1'))) OR ((E3 = '1') AND (SW3 = '1'))) OR ((E4 = '1') AND (SW4 = '1'))) OR ((E5 = '1') AND (SW5 = '1'))) OR ((E6 = '1') AND (SW6 = '1'))) OR ((E7 = '1') AND (SW7 = '1'))) OR ((E8 = '1') AND (SW8 = '1')))) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Base;
                    END IF;

                    Fermee <= '1';
                WHEN OTHERS => 
                    Fermee <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
