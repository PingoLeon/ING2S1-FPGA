-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition
-- Created on Thu Nov 02 17:26:12 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY IsArrived2sec IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        E1 : IN STD_LOGIC := '0';
        E2 : IN STD_LOGIC := '0';
        E3 : IN STD_LOGIC := '0';
        E4 : IN STD_LOGIC := '0';
        E5 : IN STD_LOGIC := '0';
        E6 : IN STD_LOGIC := '0';
        E7 : IN STD_LOGIC := '0';
        E8 : IN STD_LOGIC := '0';
        CLK2 : IN STD_LOGIC := '0';
        RESETCLOCK : OUT STD_LOGIC;
        SEC : OUT STD_LOGIC
    );
END IsArrived2sec;

ARCHITECTURE BEHAVIOR OF IsArrived2sec IS
    TYPE type_fstate IS (state4,state2,state3,state1,state6,state8,state7,state5,state15,state9);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_RESETCLOCK : STD_LOGIC := '0';
    SIGNAL reg_SEC : STD_LOGIC := '0';
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,E1,E2,E3,E4,E5,E6,E7,E8,CLK2,reg_RESETCLOCK,reg_SEC)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            reg_RESETCLOCK <= '0';
            reg_SEC <= '0';
            RESETCLOCK <= '0';
            SEC <= '0';
        ELSE
            reg_RESETCLOCK <= '0';
            reg_SEC <= '0';
            RESETCLOCK <= '0';
            SEC <= '0';
            CASE fstate IS
                WHEN state4 =>
                    IF ((CLK2 = '1')) THEN
                        reg_fstate <= state15;
                    ELSIF ((NOT((E3 = '1')) AND NOT((CLK2 = '1')))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state4;
                    END IF;

                    reg_RESETCLOCK <= '0';

                    reg_SEC <= '0';
                WHEN state2 =>
                    IF ((CLK2 = '1')) THEN
                        reg_fstate <= state15;
                    ELSIF ((NOT((E1 = '1')) AND NOT((CLK2 = '1')))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    reg_RESETCLOCK <= '0';

                    reg_SEC <= '0';
                WHEN state3 =>
                    IF ((CLK2 = '1')) THEN
                        reg_fstate <= state15;
                    ELSIF ((NOT((E2 = '1')) AND NOT((CLK2 = '1')))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    reg_RESETCLOCK <= '0';

                    reg_SEC <= '0';
                WHEN state1 =>
                    IF (((E2 = '1') AND NOT((((((((E1 = '1') OR (E3 = '1')) OR (E4 = '1')) OR (E5 = '1')) OR (E6 = '1')) OR (E7 = '1')) OR (E8 = '1'))))) THEN
                        reg_fstate <= state3;
                    ELSIF (((E1 = '1') AND NOT((((((((E2 = '1') OR (E3 = '1')) OR (E4 = '1')) OR (E5 = '1')) OR (E6 = '1')) OR (E7 = '1')) OR (E8 = '1'))))) THEN
                        reg_fstate <= state2;
                    ELSIF (((E3 = '1') AND NOT((((((((E2 = '1') OR (E1 = '1')) OR (E4 = '1')) OR (E5 = '1')) OR (E6 = '1')) OR (E7 = '1')) OR (E8 = '1'))))) THEN
                        reg_fstate <= state4;
                    ELSIF (((E4 = '1') AND NOT((((((((E2 = '1') OR (E3 = '1')) OR (E1 = '1')) OR (E5 = '1')) OR (E6 = '1')) OR (E7 = '1')) OR (E8 = '1'))))) THEN
                        reg_fstate <= state5;
                    ELSIF (((E5 = '1') AND NOT((((((((E2 = '1') OR (E3 = '1')) OR (E4 = '1')) OR (E1 = '1')) OR (E6 = '1')) OR (E7 = '1')) OR (E8 = '1'))))) THEN
                        reg_fstate <= state6;
                    ELSIF (((E6 = '1') AND NOT((((((((E2 = '1') OR (E3 = '1')) OR (E4 = '1')) OR (E5 = '1')) OR (E1 = '1')) OR (E7 = '1')) OR (E8 = '1'))))) THEN
                        reg_fstate <= state7;
                    ELSIF (((E7 = '1') AND NOT((((((((E2 = '1') OR (E3 = '1')) OR (E4 = '1')) OR (E5 = '1')) OR (E6 = '1')) OR (E1 = '1')) OR (E8 = '1'))))) THEN
                        reg_fstate <= state8;
                    ELSIF (((E8 = '1') AND NOT((((((((E2 = '1') OR (E3 = '1')) OR (E4 = '1')) OR (E5 = '1')) OR (E6 = '1')) OR (E7 = '1')) OR (E1 = '1'))))) THEN
                        reg_fstate <= state9;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    reg_RESETCLOCK <= '1';

                    reg_SEC <= '0';
                WHEN state6 =>
                    IF ((CLK2 = '1')) THEN
                        reg_fstate <= state15;
                    ELSIF ((NOT((E5 = '1')) AND NOT((CLK2 = '1')))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state6;
                    END IF;

                    reg_RESETCLOCK <= '0';

                    reg_SEC <= '0';
                WHEN state8 =>
                    IF ((CLK2 = '1')) THEN
                        reg_fstate <= state15;
                    ELSIF ((NOT((E7 = '1')) AND NOT((CLK2 = '1')))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state8;
                    END IF;

                    reg_RESETCLOCK <= '0';

                    reg_SEC <= '0';
                WHEN state7 =>
                    IF ((CLK2 = '1')) THEN
                        reg_fstate <= state15;
                    ELSIF ((NOT((E6 = '1')) AND NOT((CLK2 = '1')))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state7;
                    END IF;

                    reg_RESETCLOCK <= '0';

                    reg_SEC <= '0';
                WHEN state5 =>
                    IF ((NOT((E4 = '1')) AND NOT((CLK2 = '1')))) THEN
                        reg_fstate <= state1;
                    ELSIF ((CLK2 = '1')) THEN
                        reg_fstate <= state15;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state5;
                    END IF;

                    reg_RESETCLOCK <= '0';

                    reg_SEC <= '0';
                WHEN state15 =>
                    reg_fstate <= state15;

                    reg_RESETCLOCK <= '0';

                    reg_SEC <= '1';
                WHEN state9 =>
                    IF ((NOT((E8 = '1')) AND NOT((CLK2 = '1')))) THEN
                        reg_fstate <= state1;
                    ELSIF ((CLK2 = '1')) THEN
                        reg_fstate <= state15;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state9;
                    END IF;

                    reg_RESETCLOCK <= '0';

                    reg_SEC <= '0';
                WHEN OTHERS => 
                    reg_RESETCLOCK <= 'X';
                    reg_SEC <= 'X';
                    report "Reach undefined state";
            END CASE;
            RESETCLOCK <= reg_RESETCLOCK;
            SEC <= reg_SEC;
        END IF;
    END PROCESS;
END BEHAVIOR;
