-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition
-- Created on Tue Oct 24 17:04:53 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY A2LED IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        B1 : IN STD_LOGIC := '0';
        CLK5 : IN STD_LOGIC := '0';
        LED : OUT STD_LOGIC
    );
END A2LED;

ARCHITECTURE BEHAVIOR OF A2LED IS
    TYPE type_fstate IS (base,appui1,relache1,appui2,razappui3,relache2maintenanceactive);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_LED : STD_LOGIC := '0';
BEGIN
    PROCESS (clock,reg_fstate,reg_LED)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
            LED <= reg_LED;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,B1,CLK5)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= base;
            reg_LED <= '0';
        ELSE
            reg_LED <= '0';
            CASE fstate IS
                WHEN base =>
                    IF ((B1 = '1')) THEN
                        reg_fstate <= appui1;
                    ELSIF (NOT((B1 = '1'))) THEN
                        reg_fstate <= base;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= base;
                    END IF;

                    reg_LED <= '0';
                WHEN appui1 =>
                    IF (NOT((B1 = '1'))) THEN
                        reg_fstate <= relache1;
                    ELSIF ((B1 = '1')) THEN
                        reg_fstate <= appui1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= appui1;
                    END IF;

                    reg_LED <= '0';
                WHEN relache1 =>
                    IF (((B1 = '1') AND NOT((CLK5 = '1')))) THEN
                        reg_fstate <= appui2;
                    ELSIF ((CLK5 = '1')) THEN
                        reg_fstate <= base;
                    ELSIF ((NOT((B1 = '1')) AND NOT((CLK5 = '1')))) THEN
                        reg_fstate <= relache1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= relache1;
                    END IF;

                    reg_LED <= '0';
                WHEN appui2 =>
                    IF (NOT((B1 = '1'))) THEN
                        reg_fstate <= relache2maintenanceactive;
                    ELSIF ((B1 = '1')) THEN
                        reg_fstate <= appui2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= appui2;
                    END IF;

                    reg_LED <= '0';
                WHEN razappui3 =>
                    IF (NOT((B1 = '1'))) THEN
                        reg_fstate <= base;
                    ELSIF ((B1 = '1')) THEN
                        reg_fstate <= razappui3;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= razappui3;
                    END IF;

                    reg_LED <= '1';
                WHEN relache2maintenanceactive =>
                    IF ((B1 = '1')) THEN
                        reg_fstate <= razappui3;
                    ELSIF (NOT((B1 = '1'))) THEN
                        reg_fstate <= relache2maintenanceactive;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= relache2maintenanceactive;
                    END IF;

                    reg_LED <= '1';
                WHEN OTHERS => 
                    reg_LED <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
