-- Copyright (C) 2020  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and any partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details, at
-- https://fpgasoftware.intel.com/eula.

-- Generated by Quartus Prime Version 20.1.0 Build 711 06/05/2020 SJ Lite Edition
-- Created on Thu Nov 02 12:04:10 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Buzzer IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        LED00 : IN STD_LOGIC := '0';
        LED01 : IN STD_LOGIC := '0';
        LED02 : IN STD_LOGIC := '0';
        LED03 : IN STD_LOGIC := '0';
        LED04 : IN STD_LOGIC := '0';
        LED05 : IN STD_LOGIC := '0';
        LED06 : IN STD_LOGIC := '0';
        LED07 : IN STD_LOGIC := '0';
        buzz : OUT STD_LOGIC
    );
END Buzzer;

ARCHITECTURE BEHAVIOR OF Buzzer IS
    TYPE type_fstate IS (state1,RDC,Etage2,Etage1,Prez,Etage6,Etage3,Etage4,Etage5,buzzstate);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
    SIGNAL reg_buzz : STD_LOGIC := '0';
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,LED00,LED01,LED02,LED03,LED04,LED05,LED06,LED07,reg_buzz)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            reg_buzz <= '0';
            buzz <= '0';
        ELSE
            reg_buzz <= '0';
            buzz <= '0';
            CASE fstate IS
                WHEN state1 =>
                    IF (((((((((LED00 = '1') OR (LED01 = '1')) OR (LED02 = '1')) OR (LED03 = '1')) OR (LED04 = '1')) OR (LED05 = '1')) OR (LED06 = '1')) OR (LED07 = '1'))) THEN
                        reg_fstate <= buzzstate;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    reg_buzz <= '0';
                WHEN RDC =>
                    IF (NOT((LED00 = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= RDC;
                    END IF;

                    reg_buzz <= '0';
                WHEN Etage2 =>
                    IF (NOT((LED02 = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Etage2;
                    END IF;

                    reg_buzz <= '0';
                WHEN Etage1 =>
                    IF (NOT((LED01 = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Etage1;
                    END IF;

                    reg_buzz <= '0';
                WHEN Prez =>
                    IF (NOT((LED07 = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Prez;
                    END IF;

                    reg_buzz <= '0';
                WHEN Etage6 =>
                    IF (NOT((LED06 = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Etage6;
                    END IF;

                    reg_buzz <= '0';
                WHEN Etage3 =>
                    IF (NOT((LED03 = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Etage3;
                    END IF;

                    reg_buzz <= '0';
                WHEN Etage4 =>
                    IF (NOT((LED04 = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Etage4;
                    END IF;

                    reg_buzz <= '0';
                WHEN Etage5 =>
                    IF (NOT((LED05 = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= Etage5;
                    END IF;

                    reg_buzz <= '0';
                WHEN buzzstate =>
                    IF (((LED00 = '1') AND NOT((((((((LED01 = '1') OR (LED02 = '1')) OR (LED03 = '1')) OR (LED04 = '1')) OR (LED05 = '1')) OR (LED06 = '1')) OR (LED07 = '1'))))) THEN
                        reg_fstate <= RDC;
                    ELSIF (((LED02 = '1') AND NOT((((((((LED01 = '1') OR (LED00 = '1')) OR (LED03 = '1')) OR (LED04 = '1')) OR (LED05 = '1')) OR (LED06 = '1')) OR (LED07 = '1'))))) THEN
                        reg_fstate <= Etage2;
                    ELSIF (((LED03 = '1') AND NOT((((((((LED01 = '1') OR (LED02 = '1')) OR (LED00 = '1')) OR (LED04 = '1')) OR (LED05 = '1')) OR (LED06 = '1')) OR (LED07 = '1'))))) THEN
                        reg_fstate <= Etage3;
                    ELSIF (((LED04 = '1') AND NOT((((((((LED01 = '1') OR (LED02 = '1')) OR (LED03 = '1')) OR (LED00 = '1')) OR (LED05 = '1')) OR (LED06 = '1')) OR (LED07 = '1'))))) THEN
                        reg_fstate <= Etage4;
                    ELSIF (((LED07 = '1') AND NOT((((((((LED01 = '1') OR (LED02 = '1')) OR (LED03 = '1')) OR (LED04 = '1')) OR (LED05 = '1')) OR (LED06 = '1')) OR (LED00 = '1'))))) THEN
                        reg_fstate <= Prez;
                    ELSIF (((LED06 = '1') AND NOT((((((((LED01 = '1') OR (LED02 = '1')) OR (LED03 = '1')) OR (LED04 = '1')) OR (LED05 = '1')) OR (LED00 = '1')) OR (LED07 = '1'))))) THEN
                        reg_fstate <= Etage6;
                    ELSIF (((LED05 = '1') AND NOT((((((((LED01 = '1') OR (LED02 = '1')) OR (LED03 = '1')) OR (LED04 = '1')) OR (LED00 = '1')) OR (LED06 = '1')) OR (LED07 = '1'))))) THEN
                        reg_fstate <= Etage5;
                    ELSIF (((LED01 = '1') AND NOT((((((((LED00 = '1') OR (LED02 = '1')) OR (LED03 = '1')) OR (LED04 = '1')) OR (LED05 = '1')) OR (LED06 = '1')) OR (LED07 = '1'))))) THEN
                        reg_fstate <= Etage1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= buzzstate;
                    END IF;

                    reg_buzz <= '1';
                WHEN OTHERS => 
                    reg_buzz <= 'X';
                    report "Reach undefined state";
            END CASE;
            buzz <= reg_buzz;
        END IF;
    END PROCESS;
END BEHAVIOR;
